module run (CLOCK_50,LEDG,LEDR);
input CLOCK_50;
output reg [8:0] LEDG;
output reg [17:0] LEDR;

reg []

always @(negedge CLOCK_50)
begin 
	




end
endmodule 