module LED_state
(
	input	clk,
	output reg [7:0] LEDG,
	output reg [2:0]state
);

	
	
	
endmodule
